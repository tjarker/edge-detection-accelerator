library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;


entity Selection is
    port(
        clk: in bit_t;
        reset: in bit_t;
        
    );
end entity;